library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;
  
entity Clock_Divider is
port ( 
	clk,reset: in std_logic;
	clock_out: out std_logic);
end Clock_Divider;
  
architecture bhv of Clock_Divider is
  
signal count: integer:=1;
signal tmp : std_logic := '0';
  
begin
  
--FPGA CYCLONE IV punya freq clock 50Mhz, untuk mengsinkronkan dengan komunikasi UART 9600 bits/sec,
--Kita harus membuat frekuensi clock menjadi 872.727 Hz (agar setiap 1 periode clock, mengirim 1 bit)
--50Mhz/(2.count) = 872.72727
--Count = 28645.83, dibulatkan saja menjadi 28646.

process(clk,reset)
begin
	if(reset='1') then
	count<=1;
	tmp<='0';
	elsif(clk'event and clk='1') then
	count <=count+1;
	if (count = 28646) then 
	tmp <= NOT tmp;
	count <= 1;
	end if;
end if;
clock_out <= tmp;
end process;
  
end bhv;
